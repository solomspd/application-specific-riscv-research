module XORR(input [31:0] a,b, output[31:0] o)
o = a^b;
endmodule