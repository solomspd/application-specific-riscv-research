module alu_ctrl (input [1:0]alu_op, input [6:0]func7, input [2:0]func3, output [3:0]out);



endmodule